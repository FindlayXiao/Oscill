module char_set(
	input clk,
	input rst_n,
	input [3:0] data,
	output reg [7:0] col0,
	output reg [7:0] col1,
	output reg [7:0] col2,
	output reg [7:0] col3,
	output reg [7:0] col4,
	output reg [7:0] col5,
	output reg [7:0] col6
	);

	always @(posedge clk or negedge rst_n)
		begin
			if (!rst_n)
				begin
					col0 <= 8'b0000_0000;
					col1 <= 8'b0000_0000;
					col2 <= 8'b0000_0000;
					col3 <= 8'b0000_0000;
					col4 <= 8'b0000_0000;
					col5 <= 8'b0000_0000;
					col6 <= 8'b0000_0000;
				end
			else
				begin
					case (data)
						4'd1: // "F"
							begin
								col0 <= 8'b0000_0000;
								col1 <= 8'b0111_1111;
								col2 <= 8'b0000_1001;
								col3 <= 8'b0000_1001;
								col4 <= 8'b0000_1001;
								col5 <= 8'b0000_0001;
								col6 <= 8'b0000_0000;
							end
						4'd2: // "H"
							begin
								col0 <= 8'b0000_0000;
								col1 <= 8'b0111_1111;
								col2 <= 8'b0000_1000;
								col3 <= 8'b0000_1000;
								col4 <= 8'b0000_1000;
								col5 <= 8'b0111_1111;
								col6 <= 8'b0000_0000;
							end
						4'd3: // "I"
							begin
								col0 <= 8'b0000_0000;
								col1 <= 8'b0000_0000;
								col2 <= 8'b0100_0001;
								col3 <= 8'b0111_1111;
								col4 <= 8'b0100_0001;
								col5 <= 8'b0000_0000;
								col6 <= 8'b0000_0000;
							end
					    4'd4: // "K"
							begin
								col0 <= 8'b0000_0000;
								col1 <= 8'b0111_1111;
								col2 <= 8'b0000_1000;
								col3 <= 8'b0001_0100;
								col4 <= 8'b0010_0010;
								col5 <= 8'b0100_0001;
								col6 <= 8'b0000_0000;
							end
						4'd5: // "U"
							begin
								col0 <= 8'b0000_0000;
								col1 <= 8'b0011_1111;
								col2 <= 8'b0100_0000;
								col3 <= 8'b0100_0000;
								col4 <= 8'b0100_0000;
								col5 <= 8'b0011_1111;
								col6 <= 8'b0000_0000;
							end
						4'd6: // "Q"
							begin
								col0 <= 8'b0000_0000;
								col1 <= 8'b0011_1110;
								col2 <= 8'b0100_0001;
								col3 <= 8'b0101_0001;
								col4 <= 8'b0110_0001;
								col5 <= 8'b0111_1110;
								col6 <= 8'b0000_0000;
							end
						4'd7: // "△"
							begin
								col0 <= 8'b0000_0000;
								col1 <= 8'b0111_0000;
								col2 <= 8'b0100_1100;
								col3 <= 8'b0100_0011;
								col4 <= 8'b0100_1100;
								col5 <= 8'b0111_0000;
								col6 <= 8'b0000_0000;
							end
						4'd8: // "T"
							begin
								col0 <= 8'b0000_0000;
								col1 <= 8'b0000_0001;
								col2 <= 8'b0000_0001;
								col3 <= 8'b0111_1111;
								col4 <= 8'b0000_0001;
								col5 <= 8'b0000_0001;
								col6 <= 8'b0000_0000;
							end
						4'd9: // "V"
							begin
								col0 <= 8'b0000_0000;
								col1 <= 8'b0001_1111;
								col2 <= 8'b0010_0000;
								col3 <= 8'b0100_0000;
								col4 <= 8'b0010_0000;
								col5 <= 8'b0001_1111;
								col6 <= 8'b0000_0000;
							end
						4'd10: // "X"
							begin
								col0 <= 8'b0000_0000;
								col1 <= 8'b0110_0011;
								col2 <= 8'b0001_0100;
								col3 <= 8'b0000_1000;
								col4 <= 8'b0001_0100;
								col5 <= 8'b0110_0011;
								col6 <= 8'b0000_0000;
							end
						4'd11: // "Y"
							begin
								col0 <= 8'b0000_0000;
								col1 <= 8'b0000_0011;
								col2 <= 8'b0000_0100;
								col3 <= 8'b0111_1000;
								col4 <= 8'b0000_0100;
								col5 <= 8'b0000_0011;
								col6 <= 8'b0000_0000;
							end
						4'd12: // "Z"
							begin
								col0 <= 8'b0000_0000;
								col1 <= 8'b0110_0001;
								col2 <= 8'b0101_0001;
								col3 <= 8'b0100_1001;
								col4 <= 8'b0100_0101;
								col5 <= 8'b0100_0011;
								col6 <= 8'b0000_0000;
							end
						4'd13: // " "
							begin
								col0 <= 8'b0000_0000;
								col1 <= 8'b0000_0000;
								col2 <= 8'b0000_0000;
								col3 <= 8'b0000_0000;
								col4 <= 8'b0000_0000;
								col5 <= 8'b0000_0000;
								col6 <= 8'b0000_0000;
							end
						4'd14: // ":"
							begin
								col0 <= 8'b0000_0000;
								col1 <= 8'b0000_0000;
								col2 <= 8'b0011_0110;
								col3 <= 8'b0011_0110;
								col4 <= 8'b0000_0000;
								col5 <= 8'b0000_0000;
								col6 <= 8'b0000_0000;
							end
						4'd15: // "S"
							begin
								col0 <= 8'b0000_0000;
								col1 <= 8'b0010_0110;
								col2 <= 8'b0100_1001;
								col3 <= 8'b0100_1001;
								col4 <= 8'b0100_1001;
								col5 <= 8'b0011_0010;
								col6 <= 8'b0000_0000;
							end
						default: // "*"
							begin
								col0 <= 8'b0000_0000;
								col1 <= 8'b0010_0010;
								col2 <= 8'b0001_0100;
								col3 <= 8'b0000_1000;
								col4 <= 8'b0001_0100;
								col5 <= 8'b0010_0010;
								col6 <= 8'b0000_0000;
							end
					endcase
				end
		end

endmodule